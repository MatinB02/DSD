library verilog;
use verilog.vl_types.all;
entity tb_karatsuba_multiplier is
end tb_karatsuba_multiplier;
