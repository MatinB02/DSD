library verilog;
use verilog.vl_types.all;
entity tb_pwm_ramp is
end tb_pwm_ramp;
