library verilog;
use verilog.vl_types.all;
entity manchester_carry_chain_adder_tb is
end manchester_carry_chain_adder_tb;
